`include "defines.vh"

module W(
    input[3:0] dstE
);

endmodule 
